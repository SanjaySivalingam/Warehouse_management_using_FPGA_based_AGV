module dijkstra_mod(
    input clk,
    input [7:0] src,
    input [7:0] dest,
    output reg path_ready = 0,
    output reg [95:0] path //can accompany 12 nodes including src and dest
    );
   
   
    reg [5:0] dist [0:67] ;
    reg [67:0] visited = 0 ;
    reg [6:0] parent [0:67] ;
    reg [6:0] key = 0 ;
    reg [6:0] u = 0 ;
    reg [6:0] v = 0 ;
    reg [5:0] min = 60 ;
    integer i = 0;
    integer g = 0;
    integer j = 1 ;
    reg [6:0] index_src ;
    reg [6:0] index_dest ;
    reg [7:0] value ;
    reg [6:0] index ;
    reg [7:0] temp = 0 ;
    reg [7:0] flag2 = 0 ;
    reg done = 0 ;
    reg [6:0] n_index ;
    reg [7:0] node ;
    reg [6:0] temp_index = 0 ;
    reg [6:0] flag = 0 ;
    reg [7:0] temp_node;  
    reg [5:0]graph[0:67][0:67];

initial
    begin
      {graph[0][0],graph[0][1],graph[0][2],graph[0][3],graph[0][4],graph[0][5],graph[0][6],graph[0][7],graph[0][8],graph[0][9],graph[0][10],graph[0][11],graph[0][12],graph[0][13],graph[0][14],graph[0][15],graph[0][16],graph[0][17],graph[0][18],graph[0][19],graph[0][20],graph[0][21],graph[0][22],graph[0][23],graph[0][24],graph[0][25],graph[0][26],graph[0][27],graph[0][28],graph[0][29],graph[0][30],graph[0][31],graph[0][32],graph[0][33],graph[0][34],graph[0][35],graph[0][36], graph[0][37] , graph[0][38] , graph[0][39] , graph[0][40]  , graph[0][41] , graph[0][42] , graph[0][43] , graph[0][44] , graph[0][45] , graph[0][46] , graph[0][47] , graph[0][48] , graph[0][49] , graph[0][50] , graph[0][51] , graph[0][52] , graph[0][53] , graph[0][54] , graph[0][55] , graph[0][56] , graph[0][57] , graph[0][58] , graph[0][59] , graph[0][60] , graph[0][61] , graph[0][62] , graph[0][63] , graph[0][64] , graph[0][65] , graph[0][66], graph[0][67]} = {6'd0, 6'd60 , 6'd60, 6'd60, 6'd1, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[1][0],graph[1][1],graph[1][2],graph[1][3],graph[1][4],graph[1][5],graph[1][6],graph[1][7],graph[1][8],graph[1][9],graph[1][10],graph[1][11],graph[1][12],graph[1][13],graph[1][14],graph[1][15],graph[1][16],graph[1][17],graph[1][18],graph[1][19],graph[1][20],graph[1][21],graph[1][22],graph[1][23],graph[1][24],graph[1][25],graph[1][26],graph[1][27],graph[1][28],graph[1][29],graph[1][30],graph[1][31],graph[1][32],graph[1][33],graph[1][34],graph[1][35],graph[1][36], graph[1][37] , graph[1][38] , graph[1][39] , graph[1][40]  , graph[1][41] , graph[1][42] , graph[1][43] , graph[1][44] , graph[1][45] , graph[1][46] , graph[1][47] , graph[1][48] , graph[1][49] , graph[1][50] , graph[1][51] , graph[1][52] , graph[1][53] , graph[1][54] , graph[1][55] , graph[1][56] , graph[1][57] , graph[1][58] , graph[1][59] , graph[1][60] , graph[1][61] , graph[1][62] , graph[1][63] , graph[1][64] , graph[1][65] , graph[1][66], graph[1][67]} = {6'd60, 6'd0 , 6'd60, 6'd60, 6'd60, 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[2][0],graph[2][1],graph[2][2],graph[2][3],graph[2][4],graph[2][5],graph[2][6],graph[2][7],graph[2][8],graph[2][9],graph[2][10],graph[2][11],graph[2][12],graph[2][13],graph[2][14],graph[2][15],graph[2][16],graph[2][17],graph[2][18],graph[2][19],graph[2][20],graph[2][21],graph[2][22],graph[2][23],graph[2][24],graph[2][25],graph[2][26],graph[2][27],graph[2][28],graph[2][29],graph[2][30],graph[2][31],graph[2][32],graph[2][33],graph[2][34],graph[2][35],graph[2][36], graph[2][37] , graph[2][38] , graph[2][39] , graph[2][40]  , graph[2][41] , graph[2][42] , graph[2][43] , graph[2][44] , graph[2][45] , graph[2][46] , graph[2][47] , graph[2][48] , graph[2][49] , graph[2][50] , graph[2][51] , graph[2][52] , graph[2][53] , graph[2][54] , graph[2][55] , graph[2][56] , graph[2][57] , graph[2][58] , graph[2][59] , graph[2][60] , graph[2][61] , graph[2][62] , graph[2][63] , graph[2][64] , graph[2][65] , graph[2][66], graph[2][67]} = {6'd60, 6'd60 , 6'd0, 6'd60, 6'd60, 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[3][0],graph[3][1],graph[3][2],graph[3][3],graph[3][4],graph[3][5],graph[3][6],graph[3][7],graph[3][8],graph[3][9],graph[3][10],graph[3][11],graph[3][12],graph[3][13],graph[3][14],graph[3][15],graph[3][16],graph[3][17],graph[3][18],graph[3][19],graph[3][20],graph[3][21],graph[3][22],graph[3][23],graph[3][24],graph[3][25],graph[3][26],graph[3][27],graph[3][28],graph[3][29],graph[3][30],graph[3][31],graph[3][32],graph[3][33],graph[3][34],graph[3][35],graph[3][36], graph[3][37] , graph[3][38] , graph[3][39] , graph[3][40]  , graph[3][41] , graph[3][42] , graph[3][43] , graph[3][44] , graph[3][45] , graph[3][46] , graph[3][47] , graph[3][48] , graph[3][49] , graph[3][50] , graph[3][51] , graph[3][52] , graph[3][53] , graph[3][54] , graph[3][55] , graph[3][56] , graph[3][57] , graph[3][58] , graph[3][59] , graph[3][60] , graph[3][61] , graph[3][62] , graph[3][63] , graph[3][64] , graph[3][65] , graph[3][66], graph[3][67]} = {6'd60, 6'd60 , 6'd60, 6'd0, 6'd5, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd2 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[4][0],graph[4][1],graph[4][2],graph[4][3],graph[4][4],graph[4][5],graph[4][6],graph[4][7],graph[4][8],graph[4][9],graph[4][10],graph[4][11],graph[4][12],graph[4][13],graph[4][14],graph[4][15],graph[4][16],graph[4][17],graph[4][18],graph[4][19],graph[4][20],graph[4][21],graph[4][22],graph[4][23],graph[4][24],graph[4][25],graph[4][26],graph[4][27],graph[4][28],graph[4][29],graph[4][30],graph[4][31],graph[4][32],graph[4][33],graph[4][34],graph[4][35],graph[4][36], graph[4][37] , graph[4][38] , graph[4][39] , graph[4][40]  , graph[4][41] , graph[4][42] , graph[4][43] , graph[4][44] , graph[4][45] , graph[4][46] , graph[4][47] , graph[4][48] , graph[4][49] , graph[4][50] , graph[4][51] , graph[4][52] , graph[4][53] , graph[4][54] , graph[4][55] , graph[4][56] , graph[4][57] , graph[4][58] , graph[4][59] , graph[4][60] , graph[4][61] , graph[4][62] , graph[4][63] , graph[4][64] , graph[4][65] , graph[4][66], graph[4][67]} = {6'd1, 6'd60 , 6'd60, 6'd5, 6'd0, 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[5][0],graph[5][1],graph[5][2],graph[5][3],graph[5][4],graph[5][5],graph[5][6],graph[5][7],graph[5][8],graph[5][9],graph[5][10],graph[5][11],graph[5][12],graph[5][13],graph[5][14],graph[5][15],graph[5][16],graph[5][17],graph[5][18],graph[5][19],graph[5][20],graph[5][21],graph[5][22],graph[5][23],graph[5][24],graph[5][25],graph[5][26],graph[5][27],graph[5][28],graph[5][29],graph[5][30],graph[5][31],graph[5][32],graph[5][33],graph[5][34],graph[5][35],graph[5][36], graph[5][37] , graph[5][38] , graph[5][39] , graph[5][40]  , graph[5][41] , graph[5][42] , graph[5][43] , graph[5][44] , graph[5][45] , graph[5][46] , graph[5][47] , graph[5][48] , graph[5][49] , graph[5][50] , graph[5][51] , graph[5][52] , graph[5][53] , graph[5][54] , graph[5][55] , graph[5][56] , graph[5][57] , graph[5][58] , graph[5][59] , graph[5][60] , graph[5][61] , graph[5][62] , graph[5][63] , graph[5][64] , graph[5][65] , graph[5][66], graph[5][67]} = {6'd60, 6'd1 , 6'd60, 6'd60, 6'd1, 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[6][0],graph[6][1],graph[6][2],graph[6][3],graph[6][4],graph[6][5],graph[6][6],graph[6][7],graph[6][8],graph[6][9],graph[6][10],graph[6][11],graph[6][12],graph[6][13],graph[6][14],graph[6][15],graph[6][16],graph[6][17],graph[6][18],graph[6][19],graph[6][20],graph[6][21],graph[6][22],graph[6][23],graph[6][24],graph[6][25],graph[6][26],graph[6][27],graph[6][28],graph[6][29],graph[6][30],graph[6][31],graph[6][32],graph[6][33],graph[6][34],graph[6][35],graph[6][36], graph[6][37] , graph[6][38] , graph[6][39] , graph[6][40]  , graph[6][41] , graph[6][42] , graph[6][43] , graph[6][44] , graph[6][45] , graph[6][46] , graph[6][47] , graph[6][48] , graph[6][49] , graph[6][50] , graph[6][51] , graph[6][52] , graph[6][53] , graph[6][54] , graph[6][55] , graph[6][56] , graph[6][57] , graph[6][58] , graph[6][59] , graph[6][60] , graph[6][61] , graph[6][62] , graph[6][63] , graph[6][64] , graph[6][65] , graph[6][66], graph[6][67]} = {6'd60, 6'd60 , 6'd1, 6'd60, 6'd60, 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[7][0],graph[7][1],graph[7][2],graph[7][3],graph[7][4],graph[7][5],graph[7][6],graph[7][7],graph[7][8],graph[7][9],graph[7][10],graph[7][11],graph[7][12],graph[7][13],graph[7][14],graph[7][15],graph[7][16],graph[7][17],graph[7][18],graph[7][19],graph[7][20],graph[7][21],graph[7][22],graph[7][23],graph[7][24],graph[7][25],graph[7][26],graph[7][27],graph[7][28],graph[7][29],graph[7][30],graph[7][31],graph[7][32],graph[7][33],graph[7][34],graph[7][35],graph[7][36], graph[7][37] , graph[7][38] , graph[7][39] , graph[7][40]  , graph[7][41] , graph[7][42] , graph[7][43] , graph[7][44] , graph[7][45] , graph[7][46] , graph[7][47] , graph[7][48] , graph[7][49] , graph[7][50] , graph[7][51] , graph[7][52] , graph[7][53] , graph[7][54] , graph[7][55] , graph[7][56] , graph[7][57] , graph[7][58] , graph[7][59] , graph[7][60] , graph[7][61] , graph[7][62] , graph[7][63] , graph[7][64] , graph[7][65] , graph[7][66], graph[7][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd1 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd5 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[8][0],graph[8][1],graph[8][2],graph[8][3],graph[8][4],graph[8][5],graph[8][6],graph[8][7],graph[8][8],graph[8][9],graph[8][10],graph[8][11],graph[8][12],graph[8][13],graph[8][14],graph[8][15],graph[8][16],graph[8][17],graph[8][18],graph[8][19],graph[8][20],graph[8][21],graph[8][22],graph[8][23],graph[8][24],graph[8][25],graph[8][26],graph[8][27],graph[8][28],graph[8][29],graph[8][30],graph[8][31],graph[8][32],graph[8][33],graph[8][34],graph[8][35],graph[8][36], graph[8][37] , graph[8][38] , graph[8][39] , graph[8][40]  , graph[8][41] , graph[8][42] , graph[8][43] , graph[8][44] , graph[8][45] , graph[8][46] , graph[8][47] , graph[8][48] , graph[8][49] , graph[8][50] , graph[8][51] , graph[8][52] , graph[8][53] , graph[8][54] , graph[8][55] , graph[8][56] , graph[8][57] , graph[8][58] , graph[8][59] , graph[8][60] , graph[8][61] , graph[8][62] , graph[8][63] , graph[8][64] , graph[8][65] , graph[8][66], graph[8][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[9][0],graph[9][1],graph[9][2],graph[9][3],graph[9][4],graph[9][5],graph[9][6],graph[9][7],graph[9][8],graph[9][9],graph[9][10],graph[9][11],graph[9][12],graph[9][13],graph[9][14],graph[9][15],graph[9][16],graph[9][17],graph[9][18],graph[9][19],graph[9][20],graph[9][21],graph[9][22],graph[9][23],graph[9][24],graph[9][25],graph[9][26],graph[9][27],graph[9][28],graph[9][29],graph[9][30],graph[9][31],graph[9][32],graph[9][33],graph[9][34],graph[9][35],graph[9][36], graph[9][37] , graph[9][38] , graph[9][39] , graph[9][40]  , graph[9][41] , graph[9][42] , graph[9][43] , graph[9][44] , graph[9][45] , graph[9][46] , graph[9][47] , graph[9][48] , graph[9][49] , graph[9][50] , graph[9][51] , graph[9][52] , graph[9][53] , graph[9][54] , graph[9][55] , graph[9][56] , graph[9][57] , graph[9][58] , graph[9][59] , graph[9][60] , graph[9][61] , graph[9][62] , graph[9][63] , graph[9][64] , graph[9][65] , graph[9][66], graph[9][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[10][0],graph[10][1],graph[10][2],graph[10][3],graph[10][4],graph[10][5],graph[10][6],graph[10][7],graph[10][8],graph[10][9],graph[10][10],graph[10][11],graph[10][12],graph[10][13],graph[10][14],graph[10][15],graph[10][16],graph[10][17],graph[10][18],graph[10][19],graph[10][20],graph[10][21],graph[10][22],graph[10][23],graph[10][24],graph[10][25],graph[10][26],graph[10][27],graph[10][28],graph[10][29],graph[10][30],graph[10][31],graph[10][32],graph[10][33],graph[10][34],graph[10][35],graph[10][36], graph[10][37] , graph[10][38] , graph[10][39] , graph[10][40]  , graph[10][41] , graph[10][42] , graph[10][43] , graph[10][44] , graph[10][45] , graph[10][46] , graph[10][47] , graph[10][48] , graph[10][49] , graph[10][50] , graph[10][51] , graph[10][52] , graph[10][53] , graph[10][54] , graph[10][55] , graph[10][56] , graph[10][57] , graph[10][58] , graph[10][59] , graph[10][60] , graph[10][61] , graph[10][62] , graph[10][63] , graph[10][64] , graph[10][65] , graph[10][66], graph[10][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[11][0],graph[11][1],graph[11][2],graph[11][3],graph[11][4],graph[11][5],graph[11][6],graph[11][7],graph[11][8],graph[11][9],graph[11][10],graph[11][11],graph[11][12],graph[11][13],graph[11][14],graph[11][15],graph[11][16],graph[11][17],graph[11][18],graph[11][19],graph[11][20],graph[11][21],graph[11][22],graph[11][23],graph[11][24],graph[11][25],graph[11][26],graph[11][27],graph[11][28],graph[11][29],graph[11][30],graph[11][31],graph[11][32],graph[11][33],graph[11][34],graph[11][35],graph[11][36], graph[11][37] , graph[11][38] , graph[11][39] , graph[11][40]  , graph[11][41] , graph[11][42] , graph[11][43] , graph[11][44] , graph[11][45] , graph[11][46] , graph[11][47] , graph[11][48] , graph[11][49] , graph[11][50] , graph[11][51] , graph[11][52] , graph[11][53] , graph[11][54] , graph[11][55] , graph[11][56] , graph[11][57] , graph[11][58] , graph[11][59] , graph[11][60] , graph[11][61] , graph[11][62] , graph[11][63] , graph[11][64] , graph[11][65] , graph[11][66], graph[11][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd1, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[12][0],graph[12][1],graph[12][2],graph[12][3],graph[12][4],graph[12][5],graph[12][6],graph[12][7],graph[12][8],graph[12][9],graph[12][10],graph[12][11],graph[12][12],graph[12][13],graph[12][14],graph[12][15],graph[12][16],graph[12][17],graph[12][18],graph[12][19],graph[12][20],graph[12][21],graph[12][22],graph[12][23],graph[12][24],graph[12][25],graph[12][26],graph[12][27],graph[12][28],graph[12][29],graph[12][30],graph[12][31],graph[12][32],graph[12][33],graph[12][34],graph[12][35],graph[12][36], graph[12][37] , graph[12][38] , graph[12][39] , graph[12][40]  , graph[12][41] , graph[12][42] , graph[12][43] , graph[12][44] , graph[12][45] , graph[12][46] , graph[12][47] , graph[12][48] , graph[12][49] , graph[12][50] , graph[12][51] , graph[12][52] , graph[12][53] , graph[12][54] , graph[12][55] , graph[12][56] , graph[12][57] , graph[12][58] , graph[12][59] , graph[12][60] , graph[12][61] , graph[12][62] , graph[12][63] , graph[12][64] , graph[12][65] , graph[12][66], graph[12][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[13][0],graph[13][1],graph[13][2],graph[13][3],graph[13][4],graph[13][5],graph[13][6],graph[13][7],graph[13][8],graph[13][9],graph[13][10],graph[13][11],graph[13][12],graph[13][13],graph[13][14],graph[13][15],graph[13][16],graph[13][17],graph[13][18],graph[13][19],graph[13][20],graph[13][21],graph[13][22],graph[13][23],graph[13][24],graph[13][25],graph[13][26],graph[13][27],graph[13][28],graph[13][29],graph[13][30],graph[13][31],graph[13][32],graph[13][33],graph[13][34],graph[13][35],graph[13][36], graph[13][37] , graph[13][38] , graph[13][39] , graph[13][40]  , graph[13][41] , graph[13][42] , graph[13][43] , graph[13][44] , graph[13][45] , graph[13][46] , graph[13][47] , graph[13][48] , graph[13][49] , graph[13][50] , graph[13][51] , graph[13][52] , graph[13][53] , graph[13][54] , graph[13][55] , graph[13][56] , graph[13][57] , graph[13][58] , graph[13][59] , graph[13][60] , graph[13][61] , graph[13][62] , graph[13][63] , graph[13][64] , graph[13][65] , graph[13][66], graph[13][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[14][0],graph[14][1],graph[14][2],graph[14][3],graph[14][4],graph[14][5],graph[14][6],graph[14][7],graph[14][8],graph[14][9],graph[14][10],graph[14][11],graph[14][12],graph[14][13],graph[14][14],graph[14][15],graph[14][16],graph[14][17],graph[14][18],graph[14][19],graph[14][20],graph[14][21],graph[14][22],graph[14][23],graph[14][24],graph[14][25],graph[14][26],graph[14][27],graph[14][28],graph[14][29],graph[14][30],graph[14][31],graph[14][32],graph[14][33],graph[14][34],graph[14][35],graph[14][36], graph[14][37] , graph[14][38] , graph[14][39] , graph[14][40]  , graph[14][41] , graph[14][42] , graph[14][43] , graph[14][44] , graph[14][45] , graph[14][46] , graph[14][47] , graph[14][48] , graph[14][49] , graph[14][50] , graph[14][51] , graph[14][52] , graph[14][53] , graph[14][54] , graph[14][55] , graph[14][56] , graph[14][57] , graph[14][58] , graph[14][59] , graph[14][60] , graph[14][61] , graph[14][62] , graph[14][63] , graph[14][64] , graph[14][65] , graph[14][66], graph[14][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[15][0],graph[15][1],graph[15][2],graph[15][3],graph[15][4],graph[15][5],graph[15][6],graph[15][7],graph[15][8],graph[15][9],graph[15][10],graph[15][11],graph[15][12],graph[15][13],graph[15][14],graph[15][15],graph[15][16],graph[15][17],graph[15][18],graph[15][19],graph[15][20],graph[15][21],graph[15][22],graph[15][23],graph[15][24],graph[15][25],graph[15][26],graph[15][27],graph[15][28],graph[15][29],graph[15][30],graph[15][31],graph[15][32],graph[15][33],graph[15][34],graph[15][35],graph[15][36], graph[15][37] , graph[15][38] , graph[15][39] , graph[15][40]  , graph[15][41] , graph[15][42] , graph[15][43] , graph[15][44] , graph[15][45] , graph[15][46] , graph[15][47] , graph[15][48] , graph[15][49] , graph[15][50] , graph[15][51] , graph[15][52] , graph[15][53] , graph[15][54] , graph[15][55] , graph[15][56] , graph[15][57] , graph[15][58] , graph[15][59] , graph[15][60] , graph[15][61] , graph[15][62] , graph[15][63] , graph[15][64] , graph[15][65] , graph[15][66], graph[15][67]} = {6'd60, 6'd60 , 6'd60, 6'd2, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[16][0],graph[16][1],graph[16][2],graph[16][3],graph[16][4],graph[16][5],graph[16][6],graph[16][7],graph[16][8],graph[16][9],graph[16][10],graph[16][11],graph[16][12],graph[16][13],graph[16][14],graph[16][15],graph[16][16],graph[16][17],graph[16][18],graph[16][19],graph[16][20],graph[16][21],graph[16][22],graph[16][23],graph[16][24],graph[16][25],graph[16][26],graph[16][27],graph[16][28],graph[16][29],graph[16][30],graph[16][31],graph[16][32],graph[16][33],graph[16][34],graph[16][35],graph[16][36], graph[16][37] , graph[16][38] , graph[16][39] , graph[16][40]  , graph[16][41] , graph[16][42] , graph[16][43] , graph[16][44] , graph[16][45] , graph[16][46] , graph[16][47] , graph[16][48] , graph[16][49] , graph[16][50] , graph[16][51] , graph[16][52] , graph[16][53] , graph[16][54] , graph[16][55] , graph[16][56] , graph[16][57] , graph[16][58] , graph[16][59] , graph[16][60] , graph[16][61] , graph[16][62] , graph[16][63] , graph[16][64] , graph[16][65] , graph[16][66], graph[16][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[17][0],graph[17][1],graph[17][2],graph[17][3],graph[17][4],graph[17][5],graph[17][6],graph[17][7],graph[17][8],graph[17][9],graph[17][10],graph[17][11],graph[17][12],graph[17][13],graph[17][14],graph[17][15],graph[17][16],graph[17][17],graph[17][18],graph[17][19],graph[17][20],graph[17][21],graph[17][22],graph[17][23],graph[17][24],graph[17][25],graph[17][26],graph[17][27],graph[17][28],graph[17][29],graph[17][30],graph[17][31],graph[17][32],graph[17][33],graph[17][34],graph[17][35],graph[17][36], graph[17][37] , graph[17][38] , graph[17][39] , graph[17][40]  , graph[17][41] , graph[17][42] , graph[17][43] , graph[17][44] , graph[17][45] , graph[17][46] , graph[17][47] , graph[17][48] , graph[17][49] , graph[17][50] , graph[17][51] , graph[17][52] , graph[17][53] , graph[17][54] , graph[17][55] , graph[17][56] , graph[17][57] , graph[17][58] , graph[17][59] , graph[17][60] , graph[17][61] , graph[17][62] , graph[17][63] , graph[17][64] , graph[17][65] , graph[17][66], graph[17][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[18][0],graph[18][1],graph[18][2],graph[18][3],graph[18][4],graph[18][5],graph[18][6],graph[18][7],graph[18][8],graph[18][9],graph[18][10],graph[18][11],graph[18][12],graph[18][13],graph[18][14],graph[18][15],graph[18][16],graph[18][17],graph[18][18],graph[18][19],graph[18][20],graph[18][21],graph[18][22],graph[18][23],graph[18][24],graph[18][25],graph[18][26],graph[18][27],graph[18][28],graph[18][29],graph[18][30],graph[18][31],graph[18][32],graph[18][33],graph[18][34],graph[18][35],graph[18][36], graph[18][37] , graph[18][38] , graph[18][39] , graph[18][40]  , graph[18][41] , graph[18][42] , graph[18][43] , graph[18][44] , graph[18][45] , graph[18][46] , graph[18][47] , graph[18][48] , graph[18][49] , graph[18][50] , graph[18][51] , graph[18][52] , graph[18][53] , graph[18][54] , graph[18][55] , graph[18][56] , graph[18][57] , graph[18][58] , graph[18][59] , graph[18][60] , graph[18][61] , graph[18][62] , graph[18][63] , graph[18][64] , graph[18][65] , graph[18][66], graph[18][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[19][0],graph[19][1],graph[19][2],graph[19][3],graph[19][4],graph[19][5],graph[19][6],graph[19][7],graph[19][8],graph[19][9],graph[19][10],graph[19][11],graph[19][12],graph[19][13],graph[19][14],graph[19][15],graph[19][16],graph[19][17],graph[19][18],graph[19][19],graph[19][20],graph[19][21],graph[19][22],graph[19][23],graph[19][24],graph[19][25],graph[19][26],graph[19][27],graph[19][28],graph[19][29],graph[19][30],graph[19][31],graph[19][32],graph[19][33],graph[19][34],graph[19][35],graph[19][36], graph[19][37] , graph[19][38] , graph[19][39] , graph[19][40]  , graph[19][41] , graph[19][42] , graph[19][43] , graph[19][44] , graph[19][45] , graph[19][46] , graph[19][47] , graph[19][48] , graph[19][49] , graph[19][50] , graph[19][51] , graph[19][52] , graph[19][53] , graph[19][54] , graph[19][55] , graph[19][56] , graph[19][57] , graph[19][58] , graph[19][59] , graph[19][60] , graph[19][61] , graph[19][62] , graph[19][63] , graph[19][64] , graph[19][65] , graph[19][66], graph[19][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[20][0],graph[20][1],graph[20][2],graph[20][3],graph[20][4],graph[20][5],graph[20][6],graph[20][7],graph[20][8],graph[20][9],graph[20][10],graph[20][11],graph[20][12],graph[20][13],graph[20][14],graph[20][15],graph[20][16],graph[20][17],graph[20][18],graph[20][19],graph[20][20],graph[20][21],graph[20][22],graph[20][23],graph[20][24],graph[20][25],graph[20][26],graph[20][27],graph[20][28],graph[20][29],graph[20][30],graph[20][31],graph[20][32],graph[20][33],graph[20][34],graph[20][35],graph[20][36], graph[20][37] , graph[20][38] , graph[20][39] , graph[20][40]  , graph[20][41] , graph[20][42] , graph[20][43] , graph[20][44] , graph[20][45] , graph[20][46] , graph[20][47] , graph[20][48] , graph[20][49] , graph[20][50] , graph[20][51] , graph[20][52] , graph[20][53] , graph[20][54] , graph[20][55] , graph[20][56] , graph[20][57] , graph[20][58] , graph[20][59] , graph[20][60] , graph[20][61] , graph[20][62] , graph[20][63] , graph[20][64] , graph[20][65] , graph[20][66], graph[20][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[21][0],graph[21][1],graph[21][2],graph[21][3],graph[21][4],graph[21][5],graph[21][6],graph[21][7],graph[21][8],graph[21][9],graph[21][10],graph[21][11],graph[21][12],graph[21][13],graph[21][14],graph[21][15],graph[21][16],graph[21][17],graph[21][18],graph[21][19],graph[21][20],graph[21][21],graph[21][22],graph[21][23],graph[21][24],graph[21][25],graph[21][26],graph[21][27],graph[21][28],graph[21][29],graph[21][30],graph[21][31],graph[21][32],graph[21][33],graph[21][34],graph[21][35],graph[21][36], graph[21][37] , graph[21][38] , graph[21][39] , graph[21][40]  , graph[21][41] , graph[21][42] , graph[21][43] , graph[21][44] , graph[21][45] , graph[21][46] , graph[21][47] , graph[21][48] , graph[21][49] , graph[21][50] , graph[21][51] , graph[21][52] , graph[21][53] , graph[21][54] , graph[21][55] , graph[21][56] , graph[21][57] , graph[21][58] , graph[21][59] , graph[21][60] , graph[21][61] , graph[21][62] , graph[21][63] , graph[21][64] , graph[21][65] , graph[21][66], graph[21][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[22][0],graph[22][1],graph[22][2],graph[22][3],graph[22][4],graph[22][5],graph[22][6],graph[22][7],graph[22][8],graph[22][9],graph[22][10],graph[22][11],graph[22][12],graph[22][13],graph[22][14],graph[22][15],graph[22][16],graph[22][17],graph[22][18],graph[22][19],graph[22][20],graph[22][21],graph[22][22],graph[22][23],graph[22][24],graph[22][25],graph[22][26],graph[22][27],graph[22][28],graph[22][29],graph[22][30],graph[22][31],graph[22][32],graph[22][33],graph[22][34],graph[22][35],graph[22][36], graph[22][37] , graph[22][38] , graph[22][39] , graph[22][40]  , graph[22][41] , graph[22][42] , graph[22][43] , graph[22][44] , graph[22][45] , graph[22][46] , graph[22][47] , graph[22][48] , graph[22][49] , graph[22][50] , graph[22][51] , graph[22][52] , graph[22][53] , graph[22][54] , graph[22][55] , graph[22][56] , graph[22][57] , graph[22][58] , graph[22][59] , graph[22][60] , graph[22][61] , graph[22][62] , graph[22][63] , graph[22][64] , graph[22][65] , graph[22][66], graph[22][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[23][0],graph[23][1],graph[23][2],graph[23][3],graph[23][4],graph[23][5],graph[23][6],graph[23][7],graph[23][8],graph[23][9],graph[23][10],graph[23][11],graph[23][12],graph[23][13],graph[23][14],graph[23][15],graph[23][16],graph[23][17],graph[23][18],graph[23][19],graph[23][20],graph[23][21],graph[23][22],graph[23][23],graph[23][24],graph[23][25],graph[23][26],graph[23][27],graph[23][28],graph[23][29],graph[23][30],graph[23][31],graph[23][32],graph[23][33],graph[23][34],graph[23][35],graph[23][36], graph[23][37] , graph[23][38] , graph[23][39] , graph[23][40]  , graph[23][41] , graph[23][42] , graph[23][43] , graph[23][44] , graph[23][45] , graph[23][46] , graph[23][47] , graph[23][48] , graph[23][49] , graph[23][50] , graph[23][51] , graph[23][52] , graph[23][53] , graph[23][54] , graph[23][55] , graph[23][56] , graph[23][57] , graph[23][58] , graph[23][59] , graph[23][60] , graph[23][61] , graph[23][62] , graph[23][63] , graph[23][64] , graph[23][65] , graph[23][66], graph[23][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[24][0],graph[24][1],graph[24][2],graph[24][3],graph[24][4],graph[24][5],graph[24][6],graph[24][7],graph[24][8],graph[24][9],graph[24][10],graph[24][11],graph[24][12],graph[24][13],graph[24][14],graph[24][15],graph[24][16],graph[24][17],graph[24][18],graph[24][19],graph[24][20],graph[24][21],graph[24][22],graph[24][23],graph[24][24],graph[24][25],graph[24][26],graph[24][27],graph[24][28],graph[24][29],graph[24][30],graph[24][31],graph[24][32],graph[24][33],graph[24][34],graph[24][35],graph[24][36], graph[24][37] , graph[24][38] , graph[24][39] , graph[24][40]  , graph[24][41] , graph[24][42] , graph[24][43] , graph[24][44] , graph[24][45] , graph[24][46] , graph[24][47] , graph[24][48] , graph[24][49] , graph[24][50] , graph[24][51] , graph[24][52] , graph[24][53] , graph[24][54] , graph[24][55] , graph[24][56] , graph[24][57] , graph[24][58] , graph[24][59] , graph[24][60] , graph[24][61] , graph[24][62] , graph[24][63] , graph[24][64] , graph[24][65] , graph[24][66], graph[24][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[25][0],graph[25][1],graph[25][2],graph[25][3],graph[25][4],graph[25][5],graph[25][6],graph[25][7],graph[25][8],graph[25][9],graph[25][10],graph[25][11],graph[25][12],graph[25][13],graph[25][14],graph[25][15],graph[25][16],graph[25][17],graph[25][18],graph[25][19],graph[25][20],graph[25][21],graph[25][22],graph[25][23],graph[25][24],graph[25][25],graph[25][26],graph[25][27],graph[25][28],graph[25][29],graph[25][30],graph[25][31],graph[25][32],graph[25][33],graph[25][34],graph[25][35],graph[25][36], graph[25][37] , graph[25][38] , graph[25][39] , graph[25][40]  , graph[25][41] , graph[25][42] , graph[25][43] , graph[25][44] , graph[25][45] , graph[25][46] , graph[25][47] , graph[25][48] , graph[25][49] , graph[25][50] , graph[25][51] , graph[25][52] , graph[25][53] , graph[25][54] , graph[25][55] , graph[25][56] , graph[25][57] , graph[25][58] , graph[25][59] , graph[25][60] , graph[25][61] , graph[25][62] , graph[25][63] , graph[25][64] , graph[25][65] , graph[25][66], graph[25][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[26][0],graph[26][1],graph[26][2],graph[26][3],graph[26][4],graph[26][5],graph[26][6],graph[26][7],graph[26][8],graph[26][9],graph[26][10],graph[26][11],graph[26][12],graph[26][13],graph[26][14],graph[26][15],graph[26][16],graph[26][17],graph[26][18],graph[26][19],graph[26][20],graph[26][21],graph[26][22],graph[26][23],graph[26][24],graph[26][25],graph[26][26],graph[26][27],graph[26][28],graph[26][29],graph[26][30],graph[26][31],graph[26][32],graph[26][33],graph[26][34],graph[26][35],graph[26][36], graph[26][37] , graph[26][38] , graph[26][39] , graph[26][40]  , graph[26][41] , graph[26][42] , graph[26][43] , graph[26][44] , graph[26][45] , graph[26][46] , graph[26][47] , graph[26][48] , graph[26][49] , graph[26][50] , graph[26][51] , graph[26][52] , graph[26][53] , graph[26][54] , graph[26][55] , graph[26][56] , graph[26][57] , graph[26][58] , graph[26][59] , graph[26][60] , graph[26][61] , graph[26][62] , graph[26][63] , graph[26][64] , graph[26][65] , graph[26][66], graph[26][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[27][0],graph[27][1],graph[27][2],graph[27][3],graph[27][4],graph[27][5],graph[27][6],graph[27][7],graph[27][8],graph[27][9],graph[27][10],graph[27][11],graph[27][12],graph[27][13],graph[27][14],graph[27][15],graph[27][16],graph[27][17],graph[27][18],graph[27][19],graph[27][20],graph[27][21],graph[27][22],graph[27][23],graph[27][24],graph[27][25],graph[27][26],graph[27][27],graph[27][28],graph[27][29],graph[27][30],graph[27][31],graph[27][32],graph[27][33],graph[27][34],graph[27][35],graph[27][36], graph[27][37] , graph[27][38] , graph[27][39] , graph[27][40]  , graph[27][41] , graph[27][42] , graph[27][43] , graph[27][44] , graph[27][45] , graph[27][46] , graph[27][47] , graph[27][48] , graph[27][49] , graph[27][50] , graph[27][51] , graph[27][52] , graph[27][53] , graph[27][54] , graph[27][55] , graph[27][56] , graph[27][57] , graph[27][58] , graph[27][59] , graph[27][60] , graph[27][61] , graph[27][62] , graph[27][63] , graph[27][64] , graph[27][65] , graph[27][66], graph[27][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[28][0],graph[28][1],graph[28][2],graph[28][3],graph[28][4],graph[28][5],graph[28][6],graph[28][7],graph[28][8],graph[28][9],graph[28][10],graph[28][11],graph[28][12],graph[28][13],graph[28][14],graph[28][15],graph[28][16],graph[28][17],graph[28][18],graph[28][19],graph[28][20],graph[28][21],graph[28][22],graph[28][23],graph[28][24],graph[28][25],graph[28][26],graph[28][27],graph[28][28],graph[28][29],graph[28][30],graph[28][31],graph[28][32],graph[28][33],graph[28][34],graph[28][35],graph[28][36], graph[28][37] , graph[28][38] , graph[28][39] , graph[28][40]  , graph[28][41] , graph[28][42] , graph[28][43] , graph[28][44] , graph[28][45] , graph[28][46] , graph[28][47] , graph[28][48] , graph[28][49] , graph[28][50] , graph[28][51] , graph[28][52] , graph[28][53] , graph[28][54] , graph[28][55] , graph[28][56] , graph[28][57] , graph[28][58] , graph[28][59] , graph[28][60] , graph[28][61] , graph[28][62] , graph[28][63] , graph[28][64] , graph[28][65] , graph[28][66], graph[28][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[29][0],graph[29][1],graph[29][2],graph[29][3],graph[29][4],graph[29][5],graph[29][6],graph[29][7],graph[29][8],graph[29][9],graph[29][10],graph[29][11],graph[29][12],graph[29][13],graph[29][14],graph[29][15],graph[29][16],graph[29][17],graph[29][18],graph[29][19],graph[29][20],graph[29][21],graph[29][22],graph[29][23],graph[29][24],graph[29][25],graph[29][26],graph[29][27],graph[29][28],graph[29][29],graph[29][30],graph[29][31],graph[29][32],graph[29][33],graph[29][34],graph[29][35],graph[29][36], graph[29][37] , graph[29][38] , graph[29][39] , graph[29][40]  , graph[29][41] , graph[29][42] , graph[29][43] , graph[29][44] , graph[29][45] , graph[29][46] , graph[29][47] , graph[29][48] , graph[29][49] , graph[29][50] , graph[29][51] , graph[29][52] , graph[29][53] , graph[29][54] , graph[29][55] , graph[29][56] , graph[29][57] , graph[29][58] , graph[29][59] , graph[29][60] , graph[29][61] , graph[29][62] , graph[29][63] , graph[29][64] , graph[29][65] , graph[29][66], graph[29][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[30][0],graph[30][1],graph[30][2],graph[30][3],graph[30][4],graph[30][5],graph[30][6],graph[30][7],graph[30][8],graph[30][9],graph[30][10],graph[30][11],graph[30][12],graph[30][13],graph[30][14],graph[30][15],graph[30][16],graph[30][17],graph[30][18],graph[30][19],graph[30][20],graph[30][21],graph[30][22],graph[30][23],graph[30][24],graph[30][25],graph[30][26],graph[30][27],graph[30][28],graph[30][29],graph[30][30],graph[30][31],graph[30][32],graph[30][33],graph[30][34],graph[30][35],graph[30][36], graph[30][37] , graph[30][38] , graph[30][39] , graph[30][40]  , graph[30][41] , graph[30][42] , graph[30][43] , graph[30][44] , graph[30][45] , graph[30][46] , graph[30][47] , graph[30][48] , graph[30][49] , graph[30][50] , graph[30][51] , graph[30][52] , graph[30][53] , graph[30][54] , graph[30][55] , graph[30][56] , graph[30][57] , graph[30][58] , graph[30][59] , graph[30][60] , graph[30][61] , graph[30][62] , graph[30][63] , graph[30][64] , graph[30][65] , graph[30][66], graph[30][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[31][0],graph[31][1],graph[31][2],graph[31][3],graph[31][4],graph[31][5],graph[31][6],graph[31][7],graph[31][8],graph[31][9],graph[31][10],graph[31][11],graph[31][12],graph[31][13],graph[31][14],graph[31][15],graph[31][16],graph[31][17],graph[31][18],graph[31][19],graph[31][20],graph[31][21],graph[31][22],graph[31][23],graph[31][24],graph[31][25],graph[31][26],graph[31][27],graph[31][28],graph[31][29],graph[31][30],graph[31][31],graph[31][32],graph[31][33],graph[31][34],graph[31][35],graph[31][36], graph[31][37] , graph[31][38] , graph[31][39] , graph[31][40]  , graph[31][41] , graph[31][42] , graph[31][43] , graph[31][44] , graph[31][45] , graph[31][46] , graph[31][47] , graph[31][48] , graph[31][49] , graph[31][50] , graph[31][51] , graph[31][52] , graph[31][53] , graph[31][54] , graph[31][55] , graph[31][56] , graph[31][57] , graph[31][58] , graph[31][59] , graph[31][60] , graph[31][61] , graph[31][62] , graph[31][63] , graph[31][64] , graph[31][65] , graph[31][66], graph[31][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[32][0],graph[32][1],graph[32][2],graph[32][3],graph[32][4],graph[32][5],graph[32][6],graph[32][7],graph[32][8],graph[32][9],graph[32][10],graph[32][11],graph[32][12],graph[32][13],graph[32][14],graph[32][15],graph[32][16],graph[32][17],graph[32][18],graph[32][19],graph[32][20],graph[32][21],graph[32][22],graph[32][23],graph[32][24],graph[32][25],graph[32][26],graph[32][27],graph[32][28],graph[32][29],graph[32][30],graph[32][31],graph[32][32],graph[32][33],graph[32][34],graph[32][35],graph[32][36], graph[32][37] , graph[32][38] , graph[32][39] , graph[32][40]  , graph[32][41] , graph[32][42] , graph[32][43] , graph[32][44] , graph[32][45] , graph[32][46] , graph[32][47] , graph[32][48] , graph[32][49] , graph[32][50] , graph[32][51] , graph[32][52] , graph[32][53] , graph[32][54] , graph[32][55] , graph[32][56] , graph[32][57] , graph[32][58] , graph[32][59] , graph[32][60] , graph[32][61] , graph[32][62] , graph[32][63] , graph[32][64] , graph[32][65] , graph[32][66], graph[32][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[33][0],graph[33][1],graph[33][2],graph[33][3],graph[33][4],graph[33][5],graph[33][6],graph[33][7],graph[33][8],graph[33][9],graph[33][10],graph[33][11],graph[33][12],graph[33][13],graph[33][14],graph[33][15],graph[33][16],graph[33][17],graph[33][18],graph[33][19],graph[33][20],graph[33][21],graph[33][22],graph[33][23],graph[33][24],graph[33][25],graph[33][26],graph[33][27],graph[33][28],graph[33][29],graph[33][30],graph[33][31],graph[33][32],graph[33][33],graph[33][34],graph[33][35],graph[33][36], graph[33][37] , graph[33][38] , graph[33][39] , graph[33][40]  , graph[33][41] , graph[33][42] , graph[33][43] , graph[33][44] , graph[33][45] , graph[33][46] , graph[33][47] , graph[33][48] , graph[33][49] , graph[33][50] , graph[33][51] , graph[33][52] , graph[33][53] , graph[33][54] , graph[33][55] , graph[33][56] , graph[33][57] , graph[33][58] , graph[33][59] , graph[33][60] , graph[33][61] , graph[33][62] , graph[33][63] , graph[33][64] , graph[33][65] , graph[33][66], graph[33][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60, 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[34][0],graph[34][1],graph[34][2],graph[34][3],graph[34][4],graph[34][5],graph[34][6],graph[34][7],graph[34][8],graph[34][9],graph[34][10],graph[34][11],graph[34][12],graph[34][13],graph[34][14],graph[34][15],graph[34][16],graph[34][17],graph[34][18],graph[34][19],graph[34][20],graph[34][21],graph[34][22],graph[34][23],graph[34][24],graph[34][25],graph[34][26],graph[34][27],graph[34][28],graph[34][29],graph[34][30],graph[34][31],graph[34][32],graph[34][33],graph[34][34],graph[34][35],graph[34][36], graph[34][37] , graph[34][38] , graph[34][39] , graph[34][40]  , graph[34][41] , graph[34][42] , graph[34][43] , graph[34][44] , graph[34][45] , graph[34][46] , graph[34][47] , graph[34][48] , graph[34][49] , graph[34][50] , graph[34][51] , graph[34][52] , graph[34][53] , graph[34][54] , graph[34][55] , graph[34][56] , graph[34][57] , graph[34][58] , graph[34][59] , graph[34][60] , graph[34][61] , graph[34][62] , graph[34][63] , graph[34][64] , graph[34][65] , graph[34][66], graph[34][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[35][0],graph[35][1],graph[35][2],graph[35][3],graph[35][4],graph[35][5],graph[35][6],graph[35][7],graph[35][8],graph[35][9],graph[35][10],graph[35][11],graph[35][12],graph[35][13],graph[35][14],graph[35][15],graph[35][16],graph[35][17],graph[35][18],graph[35][19],graph[35][20],graph[35][21],graph[35][22],graph[35][23],graph[35][24],graph[35][25],graph[35][26],graph[35][27],graph[35][28],graph[35][29],graph[35][30],graph[35][31],graph[35][32],graph[35][33],graph[35][34],graph[35][35],graph[35][36], graph[35][37] , graph[35][38] , graph[35][39] , graph[35][40]  , graph[35][41] , graph[35][42] , graph[35][43] , graph[35][44] , graph[35][45] , graph[35][46] , graph[35][47] , graph[35][48] , graph[35][49] , graph[35][50] , graph[35][51] , graph[35][52] , graph[35][53] , graph[35][54] , graph[35][55] , graph[35][56] , graph[35][57] , graph[35][58] , graph[35][59] , graph[35][60] , graph[35][61] , graph[35][62] , graph[35][63] , graph[35][64] , graph[35][65] , graph[35][66], graph[35][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60, 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[36][0],graph[36][1],graph[36][2],graph[36][3],graph[36][4],graph[36][5],graph[36][6],graph[36][7],graph[36][8],graph[36][9],graph[36][10],graph[36][11],graph[36][12],graph[36][13],graph[36][14],graph[36][15],graph[36][16],graph[36][17],graph[36][18],graph[36][19],graph[36][20],graph[36][21],graph[36][22],graph[36][23],graph[36][24],graph[36][25],graph[36][26],graph[36][27],graph[36][28],graph[36][29],graph[36][30],graph[36][31],graph[36][32],graph[36][33],graph[36][34],graph[36][35],graph[36][36], graph[36][37] , graph[36][38] , graph[36][39] , graph[36][40]  , graph[36][41] , graph[36][42] , graph[36][43] , graph[36][44] , graph[36][45] , graph[36][46] , graph[36][47] , graph[36][48] , graph[36][49] , graph[36][50] , graph[36][51] , graph[36][52] , graph[36][53] , graph[36][54] , graph[36][55] , graph[36][56] , graph[36][57] , graph[36][58] , graph[36][59] , graph[36][60] , graph[36][61] , graph[36][62] , graph[36][63] , graph[36][64] , graph[36][65] , graph[36][66], graph[36][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60, 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[37][0],graph[37][1],graph[37][2],graph[37][3],graph[37][4],graph[37][5],graph[37][6],graph[37][7],graph[37][8],graph[37][9],graph[37][10],graph[37][11],graph[37][12],graph[37][13],graph[37][14],graph[37][15],graph[37][16],graph[37][17],graph[37][18],graph[37][19],graph[37][20],graph[37][21],graph[37][22],graph[37][23],graph[37][24],graph[37][25],graph[37][26],graph[37][27],graph[37][28],graph[37][29],graph[37][30],graph[37][31],graph[37][32],graph[37][33],graph[37][34],graph[37][35],graph[37][36], graph[37][37] , graph[37][38] , graph[37][39] , graph[37][40]  , graph[37][41] , graph[37][42] , graph[37][43] , graph[37][44] , graph[37][45] , graph[37][46] , graph[37][47] , graph[37][48] , graph[37][49] , graph[37][50] , graph[37][51] , graph[37][52] , graph[37][53] , graph[37][54] , graph[37][55] , graph[37][56] , graph[37][57] , graph[37][58] , graph[37][59] , graph[37][60] , graph[37][61] , graph[37][62] , graph[37][63] , graph[37][64] , graph[37][65] , graph[37][66], graph[37][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[38][0],graph[38][1],graph[38][2],graph[38][3],graph[38][4],graph[38][5],graph[38][6],graph[38][7],graph[38][8],graph[38][9],graph[38][10],graph[38][11],graph[38][12],graph[38][13],graph[38][14],graph[38][15],graph[38][16],graph[38][17],graph[38][18],graph[38][19],graph[38][20],graph[38][21],graph[38][22],graph[38][23],graph[38][24],graph[38][25],graph[38][26],graph[38][27],graph[38][28],graph[38][29],graph[38][30],graph[38][31],graph[38][32],graph[38][33],graph[38][34],graph[38][35],graph[38][36], graph[38][37] , graph[38][38] , graph[38][39] , graph[38][40]  , graph[38][41] , graph[38][42] , graph[38][43] , graph[38][44] , graph[38][45] , graph[38][46] , graph[38][47] , graph[38][48] , graph[38][49] , graph[38][50] , graph[38][51] , graph[38][52] , graph[38][53] , graph[38][54] , graph[38][55] , graph[38][56] , graph[38][57] , graph[38][58] , graph[38][59] , graph[38][60] , graph[38][61] , graph[38][62] , graph[38][63] , graph[38][64] , graph[38][65] , graph[38][66], graph[38][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd5 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd60 , 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd5 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[39][0],graph[39][1],graph[39][2],graph[39][3],graph[39][4],graph[39][5],graph[39][6],graph[39][7],graph[39][8],graph[39][9],graph[39][10],graph[39][11],graph[39][12],graph[39][13],graph[39][14],graph[39][15],graph[39][16],graph[39][17],graph[39][18],graph[39][19],graph[39][20],graph[39][21],graph[39][22],graph[39][23],graph[39][24],graph[39][25],graph[39][26],graph[39][27],graph[39][28],graph[39][29],graph[39][30],graph[39][31],graph[39][32],graph[39][33],graph[39][34],graph[39][35],graph[39][36], graph[39][37] , graph[39][38] , graph[39][39] , graph[39][40]  , graph[39][41] , graph[39][42] , graph[39][43] , graph[39][44] , graph[39][45] , graph[39][46] , graph[39][47] , graph[39][48] , graph[39][49] , graph[39][50] , graph[39][51] , graph[39][52] , graph[39][53] , graph[39][54] , graph[39][55] , graph[39][56] , graph[39][57] , graph[39][58] , graph[39][59] , graph[39][60] , graph[39][61] , graph[39][62] , graph[39][63] , graph[39][64] , graph[39][65] , graph[39][66], graph[39][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[40][0],graph[40][1],graph[40][2],graph[40][3],graph[40][4],graph[40][5],graph[40][6],graph[40][7],graph[40][8],graph[40][9],graph[40][10],graph[40][11],graph[40][12],graph[40][13],graph[40][14],graph[40][15],graph[40][16],graph[40][17],graph[40][18],graph[40][19],graph[40][20],graph[40][21],graph[40][22],graph[40][23],graph[40][24],graph[40][25],graph[40][26],graph[40][27],graph[40][28],graph[40][29],graph[40][30],graph[40][31],graph[40][32],graph[40][33],graph[40][34],graph[40][35],graph[40][36], graph[40][37] , graph[40][38] , graph[40][39] , graph[40][40]  , graph[40][41] , graph[40][42] , graph[40][43] , graph[40][44] , graph[40][45] , graph[40][46] , graph[40][47] , graph[40][48] , graph[40][49] , graph[40][50] , graph[40][51] , graph[40][52] , graph[40][53] , graph[40][54] , graph[40][55] , graph[40][56] , graph[40][57] , graph[40][58] , graph[40][59] , graph[40][60] , graph[40][61] , graph[40][62] , graph[40][63] , graph[40][64] , graph[40][65] , graph[40][66], graph[40][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[41][0],graph[41][1],graph[41][2],graph[41][3],graph[41][4],graph[41][5],graph[41][6],graph[41][7],graph[41][8],graph[41][9],graph[41][10],graph[41][11],graph[41][12],graph[41][13],graph[41][14],graph[41][15],graph[41][16],graph[41][17],graph[41][18],graph[41][19],graph[41][20],graph[41][21],graph[41][22],graph[41][23],graph[41][24],graph[41][25],graph[41][26],graph[41][27],graph[41][28],graph[41][29],graph[41][30],graph[41][31],graph[41][32],graph[41][33],graph[41][34],graph[41][35],graph[41][36], graph[41][37] , graph[41][38] , graph[41][39] , graph[41][40]  , graph[41][41] , graph[41][42] , graph[41][43] , graph[41][44] , graph[41][45] , graph[41][46] , graph[41][47] , graph[41][48] , graph[41][49] , graph[41][50] , graph[41][51] , graph[41][52] , graph[41][53] , graph[41][54] , graph[41][55] , graph[41][56] , graph[41][57] , graph[41][58] , graph[41][59] , graph[41][60] , graph[41][61] , graph[41][62] , graph[41][63] , graph[41][64] , graph[41][65] , graph[41][66], graph[41][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60, 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[42][0],graph[42][1],graph[42][2],graph[42][3],graph[42][4],graph[42][5],graph[42][6],graph[42][7],graph[42][8],graph[42][9],graph[42][10],graph[42][11],graph[42][12],graph[42][13],graph[42][14],graph[42][15],graph[42][16],graph[42][17],graph[42][18],graph[42][19],graph[42][20],graph[42][21],graph[42][22],graph[42][23],graph[42][24],graph[42][25],graph[42][26],graph[42][27],graph[42][28],graph[42][29],graph[42][30],graph[42][31],graph[42][32],graph[42][33],graph[42][34],graph[42][35],graph[42][36], graph[42][37] , graph[42][38] , graph[42][39] , graph[42][40]  , graph[42][41] , graph[42][42] , graph[42][43] , graph[42][44] , graph[42][45] , graph[42][46] , graph[42][47] , graph[42][48] , graph[42][49] , graph[42][50] , graph[42][51] , graph[42][52] , graph[42][53] , graph[42][54] , graph[42][55] , graph[42][56] , graph[42][57] , graph[42][58] , graph[42][59] , graph[42][60] , graph[42][61] , graph[42][62] , graph[42][63] , graph[42][64] , graph[42][65] , graph[42][66], graph[42][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60, 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60} ;
 {graph[43][0],graph[43][1],graph[43][2],graph[43][3],graph[43][4],graph[43][5],graph[43][6],graph[43][7],graph[43][8],graph[43][9],graph[43][10],graph[43][11],graph[43][12],graph[43][13],graph[43][14],graph[43][15],graph[43][16],graph[43][17],graph[43][18],graph[43][19],graph[43][20],graph[43][21],graph[43][22],graph[43][23],graph[43][24],graph[43][25],graph[43][26],graph[43][27],graph[43][28],graph[43][29],graph[43][30],graph[43][31],graph[43][32],graph[43][33],graph[43][34],graph[43][35],graph[43][36], graph[43][37] , graph[43][38] , graph[43][39] , graph[43][40]  , graph[43][41] , graph[43][42] , graph[43][43] , graph[43][44] , graph[43][45] , graph[43][46] , graph[43][47] , graph[43][48] , graph[43][49] , graph[43][50] , graph[43][51] , graph[43][52] , graph[43][53] , graph[43][54] , graph[43][55] , graph[43][56] , graph[43][57] , graph[43][58] , graph[43][59] , graph[43][60] , graph[43][61] , graph[43][62] , graph[43][63] , graph[43][64] , graph[43][65] , graph[43][66], graph[43][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[44][0],graph[44][1],graph[44][2],graph[44][3],graph[44][4],graph[44][5],graph[44][6],graph[44][7],graph[44][8],graph[44][9],graph[44][10],graph[44][11],graph[44][12],graph[44][13],graph[44][14],graph[44][15],graph[44][16],graph[44][17],graph[44][18],graph[44][19],graph[44][20],graph[44][21],graph[44][22],graph[44][23],graph[44][24],graph[44][25],graph[44][26],graph[44][27],graph[44][28],graph[44][29],graph[44][30],graph[44][31],graph[44][32],graph[44][33],graph[44][34],graph[44][35],graph[44][36], graph[44][37] , graph[44][38] , graph[44][39] , graph[44][40]  , graph[44][41] , graph[44][42] , graph[44][43] , graph[44][44] , graph[44][45] , graph[44][46] , graph[44][47] , graph[44][48] , graph[44][49] , graph[44][50] , graph[44][51] , graph[44][52] , graph[44][53] , graph[44][54] , graph[44][55] , graph[44][56] , graph[44][57] , graph[44][58] , graph[44][59] , graph[44][60] , graph[44][61] , graph[44][62] , graph[44][63] , graph[44][64] , graph[44][65] , graph[44][66], graph[44][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[45][0],graph[45][1],graph[45][2],graph[45][3],graph[45][4],graph[45][5],graph[45][6],graph[45][7],graph[45][8],graph[45][9],graph[45][10],graph[45][11],graph[45][12],graph[45][13],graph[45][14],graph[45][15],graph[45][16],graph[45][17],graph[45][18],graph[45][19],graph[45][20],graph[45][21],graph[45][22],graph[45][23],graph[45][24],graph[45][25],graph[45][26],graph[45][27],graph[45][28],graph[45][29],graph[45][30],graph[45][31],graph[45][32],graph[45][33],graph[45][34],graph[45][35],graph[45][36], graph[45][37] , graph[45][38] , graph[45][39] , graph[45][40]  , graph[45][41] , graph[45][42] , graph[45][43] , graph[45][44] , graph[45][45] , graph[45][46] , graph[45][47] , graph[45][48] , graph[45][49] , graph[45][50] , graph[45][51] , graph[45][52] , graph[45][53] , graph[45][54] , graph[45][55] , graph[45][56] , graph[45][57] , graph[45][58] , graph[45][59] , graph[45][60] , graph[45][61] , graph[45][62] , graph[45][63] , graph[45][64] , graph[45][65] , graph[45][66], graph[45][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[46][0],graph[46][1],graph[46][2],graph[46][3],graph[46][4],graph[46][5],graph[46][6],graph[46][7],graph[46][8],graph[46][9],graph[46][10],graph[46][11],graph[46][12],graph[46][13],graph[46][14],graph[46][15],graph[46][16],graph[46][17],graph[46][18],graph[46][19],graph[46][20],graph[46][21],graph[46][22],graph[46][23],graph[46][24],graph[46][25],graph[46][26],graph[46][27],graph[46][28],graph[46][29],graph[46][30],graph[46][31],graph[46][32],graph[46][33],graph[46][34],graph[46][35],graph[46][36], graph[46][37] , graph[46][38] , graph[46][39] , graph[46][40]  , graph[46][41] , graph[46][42] , graph[46][43] , graph[46][44] , graph[46][45] , graph[46][46] , graph[46][47] , graph[46][48] , graph[46][49] , graph[46][50] , graph[46][51] , graph[46][52] , graph[46][53] , graph[46][54] , graph[46][55] , graph[46][56] , graph[46][57] , graph[46][58] , graph[46][59] , graph[46][60] , graph[46][61] , graph[46][62] , graph[46][63] , graph[46][64] , graph[46][65] , graph[46][66], graph[46][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[47][0],graph[47][1],graph[47][2],graph[47][3],graph[47][4],graph[47][5],graph[47][6],graph[47][7],graph[47][8],graph[47][9],graph[47][10],graph[47][11],graph[47][12],graph[47][13],graph[47][14],graph[47][15],graph[47][16],graph[47][17],graph[47][18],graph[47][19],graph[47][20],graph[47][21],graph[47][22],graph[47][23],graph[47][24],graph[47][25],graph[47][26],graph[47][27],graph[47][28],graph[47][29],graph[47][30],graph[47][31],graph[47][32],graph[47][33],graph[47][34],graph[47][35],graph[47][36], graph[47][37] , graph[47][38] , graph[47][39] , graph[47][40]  , graph[47][41] , graph[47][42] , graph[47][43] , graph[47][44] , graph[47][45] , graph[47][46] , graph[47][47] , graph[47][48] , graph[47][49] , graph[47][50] , graph[47][51] , graph[47][52] , graph[47][53] , graph[47][54] , graph[47][55] , graph[47][56] , graph[47][57] , graph[47][58] , graph[47][59] , graph[47][60] , graph[47][61] , graph[47][62] , graph[47][63] , graph[47][64] , graph[47][65] , graph[47][66], graph[47][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[48][0],graph[48][1],graph[48][2],graph[48][3],graph[48][4],graph[48][5],graph[48][6],graph[48][7],graph[48][8],graph[48][9],graph[48][10],graph[48][11],graph[48][12],graph[48][13],graph[48][14],graph[48][15],graph[48][16],graph[48][17],graph[48][18],graph[48][19],graph[48][20],graph[48][21],graph[48][22],graph[48][23],graph[48][24],graph[48][25],graph[48][26],graph[48][27],graph[48][28],graph[48][29],graph[48][30],graph[48][31],graph[48][32],graph[48][33],graph[48][34],graph[48][35],graph[48][36], graph[48][37] , graph[48][38] , graph[48][39] , graph[48][40]  , graph[48][41] , graph[48][42] , graph[48][43] , graph[48][44] , graph[48][45] , graph[48][46] , graph[48][47] , graph[48][48] , graph[48][49] , graph[48][50] , graph[48][51] , graph[48][52] , graph[48][53] , graph[48][54] , graph[48][55] , graph[48][56] , graph[48][57] , graph[48][58] , graph[48][59] , graph[48][60] , graph[48][61] , graph[48][62] , graph[48][63] , graph[48][64] , graph[48][65] , graph[48][66], graph[48][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[49][0],graph[49][1],graph[49][2],graph[49][3],graph[49][4],graph[49][5],graph[49][6],graph[49][7],graph[49][8],graph[49][9],graph[49][10],graph[49][11],graph[49][12],graph[49][13],graph[49][14],graph[49][15],graph[49][16],graph[49][17],graph[49][18],graph[49][19],graph[49][20],graph[49][21],graph[49][22],graph[49][23],graph[49][24],graph[49][25],graph[49][26],graph[49][27],graph[49][28],graph[49][29],graph[49][30],graph[49][31],graph[49][32],graph[49][33],graph[49][34],graph[49][35],graph[49][36], graph[49][37] , graph[49][38] , graph[49][39] , graph[49][40]  , graph[49][41] , graph[49][42] , graph[49][43] , graph[49][44] , graph[49][45] , graph[49][46] , graph[49][47] , graph[49][48] , graph[49][49] , graph[49][50] , graph[49][51] , graph[49][52] , graph[49][53] , graph[49][54] , graph[49][55] , graph[49][56] , graph[49][57] , graph[49][58] , graph[49][59] , graph[49][60] , graph[49][61] , graph[49][62] , graph[49][63] , graph[49][64] , graph[49][65] , graph[49][66], graph[49][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd2 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[50][0],graph[50][1],graph[50][2],graph[50][3],graph[50][4],graph[50][5],graph[50][6],graph[50][7],graph[50][8],graph[50][9],graph[50][10],graph[50][11],graph[50][12],graph[50][13],graph[50][14],graph[50][15],graph[50][16],graph[50][17],graph[50][18],graph[50][19],graph[50][20],graph[50][21],graph[50][22],graph[50][23],graph[50][24],graph[50][25],graph[50][26],graph[50][27],graph[50][28],graph[50][29],graph[50][30],graph[50][31],graph[50][32],graph[50][33],graph[50][34],graph[50][35],graph[50][36], graph[50][37] , graph[50][38] , graph[50][39] , graph[50][40]  , graph[50][41] , graph[50][42] , graph[50][43] , graph[50][44] , graph[50][45] , graph[50][46] , graph[50][47] , graph[50][48] , graph[50][49] , graph[50][50] , graph[50][51] , graph[50][52] , graph[50][53] , graph[50][54] , graph[50][55] , graph[50][56] , graph[50][57] , graph[50][58] , graph[50][59] , graph[50][60] , graph[50][61] , graph[50][62] , graph[50][63] , graph[50][64] , graph[50][65] , graph[50][66], graph[50][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[51][0],graph[51][1],graph[51][2],graph[51][3],graph[51][4],graph[51][5],graph[51][6],graph[51][7],graph[51][8],graph[51][9],graph[51][10],graph[51][11],graph[51][12],graph[51][13],graph[51][14],graph[51][15],graph[51][16],graph[51][17],graph[51][18],graph[51][19],graph[51][20],graph[51][21],graph[51][22],graph[51][23],graph[51][24],graph[51][25],graph[51][26],graph[51][27],graph[51][28],graph[51][29],graph[51][30],graph[51][31],graph[51][32],graph[51][33],graph[51][34],graph[51][35],graph[51][36], graph[51][37] , graph[51][38] , graph[51][39] , graph[51][40]  , graph[51][41] , graph[51][42] , graph[51][43] , graph[51][44] , graph[51][45] , graph[51][46] , graph[51][47] , graph[51][48] , graph[51][49] , graph[51][50] , graph[51][51] , graph[51][52] , graph[51][53] , graph[51][54] , graph[51][55] , graph[51][56] , graph[51][57] , graph[51][58] , graph[51][59] , graph[51][60] , graph[51][61] , graph[51][62] , graph[51][63] , graph[51][64] , graph[51][65] , graph[51][66], graph[51][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[52][0],graph[52][1],graph[52][2],graph[52][3],graph[52][4],graph[52][5],graph[52][6],graph[52][7],graph[52][8],graph[52][9],graph[52][10],graph[52][11],graph[52][12],graph[52][13],graph[52][14],graph[52][15],graph[52][16],graph[52][17],graph[52][18],graph[52][19],graph[52][20],graph[52][21],graph[52][22],graph[52][23],graph[52][24],graph[52][25],graph[52][26],graph[52][27],graph[52][28],graph[52][29],graph[52][30],graph[52][31],graph[52][32],graph[52][33],graph[52][34],graph[52][35],graph[52][36], graph[52][37] , graph[52][38] , graph[52][39] , graph[52][40]  , graph[52][41] , graph[52][42] , graph[52][43] , graph[52][44] , graph[52][45] , graph[52][46] , graph[52][47] , graph[52][48] , graph[52][49] , graph[52][50] , graph[52][51] , graph[52][52] , graph[52][53] , graph[52][54] , graph[52][55] , graph[52][56] , graph[52][57] , graph[52][58] , graph[52][59] , graph[52][60] , graph[52][61] , graph[52][62] , graph[52][63] , graph[52][64] , graph[52][65] , graph[52][66], graph[52][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[53][0],graph[53][1],graph[53][2],graph[53][3],graph[53][4],graph[53][5],graph[53][6],graph[53][7],graph[53][8],graph[53][9],graph[53][10],graph[53][11],graph[53][12],graph[53][13],graph[53][14],graph[53][15],graph[53][16],graph[53][17],graph[53][18],graph[53][19],graph[53][20],graph[53][21],graph[53][22],graph[53][23],graph[53][24],graph[53][25],graph[53][26],graph[53][27],graph[53][28],graph[53][29],graph[53][30],graph[53][31],graph[53][32],graph[53][33],graph[53][34],graph[53][35],graph[53][36], graph[53][37] , graph[53][38] , graph[53][39] , graph[53][40]  , graph[53][41] , graph[53][42] , graph[53][43] , graph[53][44] , graph[53][45] , graph[53][46] , graph[53][47] , graph[53][48] , graph[53][49] , graph[53][50] , graph[53][51] , graph[53][52] , graph[53][53] , graph[53][54] , graph[53][55] , graph[53][56] , graph[53][57] , graph[53][58] , graph[53][59] , graph[53][60] , graph[53][61] , graph[53][62] , graph[53][63] , graph[53][64] , graph[53][65] , graph[53][66], graph[53][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd3 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[54][0],graph[54][1],graph[54][2],graph[54][3],graph[54][4],graph[54][5],graph[54][6],graph[54][7],graph[54][8],graph[54][9],graph[54][10],graph[54][11],graph[54][12],graph[54][13],graph[54][14],graph[54][15],graph[54][16],graph[54][17],graph[54][18],graph[54][19],graph[54][20],graph[54][21],graph[54][22],graph[54][23],graph[54][24],graph[54][25],graph[54][26],graph[54][27],graph[54][28],graph[54][29],graph[54][30],graph[54][31],graph[54][32],graph[54][33],graph[54][34],graph[54][35],graph[54][36], graph[54][37] , graph[54][38] , graph[54][39] , graph[54][40]  , graph[54][41] , graph[54][42] , graph[54][43] , graph[54][44] , graph[54][45] , graph[54][46] , graph[54][47] , graph[54][48] , graph[54][49] , graph[54][50] , graph[54][51] , graph[54][52] , graph[54][53] , graph[54][54] , graph[54][55] , graph[54][56] , graph[54][57] , graph[54][58] , graph[54][59] , graph[54][60] , graph[54][61] , graph[54][62] , graph[54][63] , graph[54][64] , graph[54][65] , graph[54][66], graph[54][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[55][0],graph[55][1],graph[55][2],graph[55][3],graph[55][4],graph[55][5],graph[55][6],graph[55][7],graph[55][8],graph[55][9],graph[55][10],graph[55][11],graph[55][12],graph[55][13],graph[55][14],graph[55][15],graph[55][16],graph[55][17],graph[55][18],graph[55][19],graph[55][20],graph[55][21],graph[55][22],graph[55][23],graph[55][24],graph[55][25],graph[55][26],graph[55][27],graph[55][28],graph[55][29],graph[55][30],graph[55][31],graph[55][32],graph[55][33],graph[55][34],graph[55][35],graph[55][36], graph[55][37] , graph[55][38] , graph[55][39] , graph[55][40]  , graph[55][41] , graph[55][42] , graph[55][43] , graph[55][44] , graph[55][45] , graph[55][46] , graph[55][47] , graph[55][48] , graph[55][49] , graph[55][50] , graph[55][51] , graph[55][52] , graph[55][53] , graph[55][54] , graph[55][55] , graph[55][56] , graph[55][57] , graph[55][58] , graph[55][59] , graph[55][60] , graph[55][61] , graph[55][62] , graph[55][63] , graph[55][64] , graph[55][65] , graph[55][66], graph[55][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[56][0],graph[56][1],graph[56][2],graph[56][3],graph[56][4],graph[56][5],graph[56][6],graph[56][7],graph[56][8],graph[56][9],graph[56][10],graph[56][11],graph[56][12],graph[56][13],graph[56][14],graph[56][15],graph[56][16],graph[56][17],graph[56][18],graph[56][19],graph[56][20],graph[56][21],graph[56][22],graph[56][23],graph[56][24],graph[56][25],graph[56][26],graph[56][27],graph[56][28],graph[56][29],graph[56][30],graph[56][31],graph[56][32],graph[56][33],graph[56][34],graph[56][35],graph[56][36], graph[56][37] , graph[56][38] , graph[56][39] , graph[56][40]  , graph[56][41] , graph[56][42] , graph[56][43] , graph[56][44] , graph[56][45] , graph[56][46] , graph[56][47] , graph[56][48] , graph[56][49] , graph[56][50] , graph[56][51] , graph[56][52] , graph[56][53] , graph[56][54] , graph[56][55] , graph[56][56] , graph[56][57] , graph[56][58] , graph[56][59] , graph[56][60] , graph[56][61] , graph[56][62] , graph[56][63] , graph[56][64] , graph[56][65] , graph[56][66], graph[56][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[57][0],graph[57][1],graph[57][2],graph[57][3],graph[57][4],graph[57][5],graph[57][6],graph[57][7],graph[57][8],graph[57][9],graph[57][10],graph[57][11],graph[57][12],graph[57][13],graph[57][14],graph[57][15],graph[57][16],graph[57][17],graph[57][18],graph[57][19],graph[57][20],graph[57][21],graph[57][22],graph[57][23],graph[57][24],graph[57][25],graph[57][26],graph[57][27],graph[57][28],graph[57][29],graph[57][30],graph[57][31],graph[57][32],graph[57][33],graph[57][34],graph[57][35],graph[57][36], graph[57][37] , graph[57][38] , graph[57][39] , graph[57][40]  , graph[57][41] , graph[57][42] , graph[57][43] , graph[57][44] , graph[57][45] , graph[57][46] , graph[57][47] , graph[57][48] , graph[57][49] , graph[57][50] , graph[57][51] , graph[57][52] , graph[57][53] , graph[57][54] , graph[57][55] , graph[57][56] , graph[57][57] , graph[57][58] , graph[57][59] , graph[57][60] , graph[57][61] , graph[57][62] , graph[57][63] , graph[57][64] , graph[57][65] , graph[57][66], graph[57][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[58][0],graph[58][1],graph[58][2],graph[58][3],graph[58][4],graph[58][5],graph[58][6],graph[58][7],graph[58][8],graph[58][9],graph[58][10],graph[58][11],graph[58][12],graph[58][13],graph[58][14],graph[58][15],graph[58][16],graph[58][17],graph[58][18],graph[58][19],graph[58][20],graph[58][21],graph[58][22],graph[58][23],graph[58][24],graph[58][25],graph[58][26],graph[58][27],graph[58][28],graph[58][29],graph[58][30],graph[58][31],graph[58][32],graph[58][33],graph[58][34],graph[58][35],graph[58][36], graph[58][37] , graph[58][38] , graph[58][39] , graph[58][40]  , graph[58][41] , graph[58][42] , graph[58][43] , graph[58][44] , graph[58][45] , graph[58][46] , graph[58][47] , graph[58][48] , graph[58][49] , graph[58][50] , graph[58][51] , graph[58][52] , graph[58][53] , graph[58][54] , graph[58][55] , graph[58][56] , graph[58][57] , graph[58][58] , graph[58][59] , graph[58][60] , graph[58][61] , graph[58][62] , graph[58][63] , graph[58][64] , graph[58][65] , graph[58][66], graph[58][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[59][0],graph[59][1],graph[59][2],graph[59][3],graph[59][4],graph[59][5],graph[59][6],graph[59][7],graph[59][8],graph[59][9],graph[59][10],graph[59][11],graph[59][12],graph[59][13],graph[59][14],graph[59][15],graph[59][16],graph[59][17],graph[59][18],graph[59][19],graph[59][20],graph[59][21],graph[59][22],graph[59][23],graph[59][24],graph[59][25],graph[59][26],graph[59][27],graph[59][28],graph[59][29],graph[59][30],graph[59][31],graph[59][32],graph[59][33],graph[59][34],graph[59][35],graph[59][36], graph[59][37] , graph[59][38] , graph[59][39] , graph[59][40]  , graph[59][41] , graph[59][42] , graph[59][43] , graph[59][44] , graph[59][45] , graph[59][46] , graph[59][47] , graph[59][48] , graph[59][49] , graph[59][50] , graph[59][51] , graph[59][52] , graph[59][53] , graph[59][54] , graph[59][55] , graph[59][56] , graph[59][57] , graph[59][58] , graph[59][59] , graph[59][60] , graph[59][61] , graph[59][62] , graph[59][63] , graph[59][64] , graph[59][65] , graph[59][66], graph[59][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[60][0],graph[60][1],graph[60][2],graph[60][3],graph[60][4],graph[60][5],graph[60][6],graph[60][7],graph[60][8],graph[60][9],graph[60][10],graph[60][11],graph[60][12],graph[60][13],graph[60][14],graph[60][15],graph[60][16],graph[60][17],graph[60][18],graph[60][19],graph[60][20],graph[60][21],graph[60][22],graph[60][23],graph[60][24],graph[60][25],graph[60][26],graph[60][27],graph[60][28],graph[60][29],graph[60][30],graph[60][31],graph[60][32],graph[60][33],graph[60][34],graph[60][35],graph[60][36], graph[60][37] , graph[60][38] , graph[60][39] , graph[60][40]  , graph[60][41] , graph[60][42] , graph[60][43] , graph[60][44] , graph[60][45] , graph[60][46] , graph[60][47] , graph[60][48] , graph[60][49] , graph[60][50] , graph[60][51] , graph[60][52] , graph[60][53] , graph[60][54] , graph[60][55] , graph[60][56] , graph[60][57] , graph[60][58] , graph[60][59] , graph[60][60] , graph[60][61] , graph[60][62] , graph[60][63] , graph[60][64] , graph[60][65] , graph[60][66], graph[60][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd2 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd5 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60};
 {graph[61][0],graph[61][1],graph[61][2],graph[61][3],graph[61][4],graph[61][5],graph[61][6],graph[61][7],graph[61][8],graph[61][9],graph[61][10],graph[61][11],graph[61][12],graph[61][13],graph[61][14],graph[61][15],graph[61][16],graph[61][17],graph[61][18],graph[61][19],graph[61][20],graph[61][21],graph[61][22],graph[61][23],graph[61][24],graph[61][25],graph[61][26],graph[61][27],graph[61][28],graph[61][29],graph[61][30],graph[61][31],graph[61][32],graph[61][33],graph[61][34],graph[61][35],graph[61][36], graph[61][37] , graph[61][38] , graph[61][39] , graph[61][40]  , graph[61][41] , graph[61][42] , graph[61][43] , graph[61][44] , graph[61][45] , graph[61][46] , graph[61][47] , graph[61][48] , graph[61][49] , graph[61][50] , graph[61][51] , graph[61][52] , graph[61][53] , graph[61][54] , graph[61][55] , graph[61][56] , graph[61][57] , graph[61][58] , graph[61][59] , graph[61][60] , graph[61][61] , graph[61][62] , graph[61][63] , graph[61][64] , graph[61][65] , graph[61][66], graph[61][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd5 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60};
 {graph[62][0],graph[62][1],graph[62][2],graph[62][3],graph[62][4],graph[62][5],graph[62][6],graph[62][7],graph[62][8],graph[62][9],graph[62][10],graph[62][11],graph[62][12],graph[62][13],graph[62][14],graph[62][15],graph[62][16],graph[62][17],graph[62][18],graph[62][19],graph[62][20],graph[62][21],graph[62][22],graph[62][23],graph[62][24],graph[62][25],graph[62][26],graph[62][27],graph[62][28],graph[62][29],graph[62][30],graph[62][31],graph[62][32],graph[62][33],graph[62][34],graph[62][35],graph[62][36], graph[62][37] , graph[62][38] , graph[62][39] , graph[62][40]  , graph[62][41] , graph[62][42] , graph[62][43] , graph[62][44] , graph[62][45] , graph[62][46] , graph[62][47] , graph[62][48] , graph[62][49] , graph[62][50] , graph[62][51] , graph[62][52] , graph[62][53] , graph[62][54] , graph[62][55] , graph[62][56] , graph[62][57] , graph[62][58] , graph[62][59] , graph[62][60] , graph[62][61] , graph[62][62] , graph[62][63] , graph[62][64] , graph[62][65] , graph[62][66], graph[62][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd60};
 {graph[63][0],graph[63][1],graph[63][2],graph[63][3],graph[63][4],graph[63][5],graph[63][6],graph[63][7],graph[63][8],graph[63][9],graph[63][10],graph[63][11],graph[63][12],graph[63][13],graph[63][14],graph[63][15],graph[63][16],graph[63][17],graph[63][18],graph[63][19],graph[63][20],graph[63][21],graph[63][22],graph[63][23],graph[63][24],graph[63][25],graph[63][26],graph[63][27],graph[63][28],graph[63][29],graph[63][30],graph[63][31],graph[63][32],graph[63][33],graph[63][34],graph[63][35],graph[63][36], graph[63][37] , graph[63][38] , graph[63][39] , graph[63][40]  , graph[63][41] , graph[63][42] , graph[63][43] , graph[63][44] , graph[63][45] , graph[63][46] , graph[63][47] , graph[63][48] , graph[63][49] , graph[63][50] , graph[63][51] , graph[63][52] , graph[63][53] , graph[63][54] , graph[63][55] , graph[63][56] , graph[63][57] , graph[63][58] , graph[63][59] , graph[63][60] , graph[63][61] , graph[63][62] , graph[63][63] , graph[63][64] , graph[63][65] , graph[63][66], graph[63][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd1 , 6'd60 , 6'd60 , 6'd1};
 {graph[64][0],graph[64][1],graph[64][2],graph[64][3],graph[64][4],graph[64][5],graph[64][6],graph[64][7],graph[64][8],graph[64][9],graph[64][10],graph[64][11],graph[64][12],graph[64][13],graph[64][14],graph[64][15],graph[64][16],graph[64][17],graph[64][18],graph[64][19],graph[64][20],graph[64][21],graph[64][22],graph[64][23],graph[64][24],graph[64][25],graph[64][26],graph[64][27],graph[64][28],graph[64][29],graph[64][30],graph[64][31],graph[64][32],graph[64][33],graph[64][34],graph[64][35],graph[64][36], graph[64][37] , graph[64][38] , graph[64][39] , graph[64][40]  , graph[64][41] , graph[64][42] , graph[64][43] , graph[64][44] , graph[64][45] , graph[64][46] , graph[64][47] , graph[64][48] , graph[64][49] , graph[64][50] , graph[64][51] , graph[64][52] , graph[64][53] , graph[64][54] , graph[64][55] , graph[64][56] , graph[64][57] , graph[64][58] , graph[64][59] , graph[64][60] , graph[64][61] , graph[64][62] , graph[64][63] , graph[64][64] , graph[64][65] , graph[64][66], graph[64][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd5 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd0 , 6'd60 , 6'd60 , 6'd60};
 {graph[65][0],graph[65][1],graph[65][2],graph[65][3],graph[65][4],graph[65][5],graph[65][6],graph[65][7],graph[65][8],graph[65][9],graph[65][10],graph[65][11],graph[65][12],graph[65][13],graph[65][14],graph[65][15],graph[65][16],graph[65][17],graph[65][18],graph[65][19],graph[65][20],graph[65][21],graph[65][22],graph[65][23],graph[65][24],graph[65][25],graph[65][26],graph[65][27],graph[65][28],graph[65][29],graph[65][30],graph[65][31],graph[65][32],graph[65][33],graph[65][34],graph[65][35],graph[65][36], graph[65][37] , graph[65][38] , graph[65][39] , graph[65][40]  , graph[65][41] , graph[65][42] , graph[65][43] , graph[65][44] , graph[65][45] , graph[65][46] , graph[65][47] , graph[65][48] , graph[65][49] , graph[65][50] , graph[65][51] , graph[65][52] , graph[65][53] , graph[65][54] , graph[65][55] , graph[65][56] , graph[65][57] , graph[65][58] , graph[65][59] , graph[65][60] , graph[65][61] , graph[65][62] , graph[65][63] , graph[65][64] , graph[65][65] , graph[65][66], graph[65][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60 , 6'd60};
 {graph[66][0],graph[66][1],graph[66][2],graph[66][3],graph[66][4],graph[66][5],graph[66][6],graph[66][7],graph[66][8],graph[66][9],graph[66][10],graph[66][11],graph[66][12],graph[66][13],graph[66][14],graph[66][15],graph[66][16],graph[66][17],graph[66][18],graph[66][19],graph[66][20],graph[66][21],graph[66][22],graph[66][23],graph[66][24],graph[66][25],graph[66][26],graph[66][27],graph[66][28],graph[66][29],graph[66][30],graph[66][31],graph[66][32],graph[66][33],graph[66][34],graph[66][35],graph[66][36], graph[66][37] , graph[66][38] , graph[66][39] , graph[66][40]  , graph[66][41] , graph[66][42] , graph[66][43] , graph[66][44] , graph[66][45] , graph[66][46] , graph[66][47] , graph[66][48] , graph[66][49] , graph[66][50] , graph[66][51] , graph[66][52] , graph[66][53] , graph[66][54] , graph[66][55] , graph[66][56] , graph[66][57] , graph[66][58] , graph[66][59] , graph[66][60] , graph[66][61] , graph[66][62] , graph[66][63] , graph[66][64] , graph[66][65] , graph[66][66], graph[66][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0 , 6'd60};
 {graph[67][0],graph[67][1],graph[67][2],graph[67][3],graph[67][4],graph[67][5],graph[67][6],graph[67][7],graph[67][8],graph[67][9],graph[67][10],graph[67][11],graph[67][12],graph[67][13],graph[67][14],graph[67][15],graph[67][16],graph[67][17],graph[67][18],graph[67][19],graph[67][20],graph[67][21],graph[67][22],graph[67][23],graph[67][24],graph[67][25],graph[67][26],graph[67][27],graph[67][28],graph[67][29],graph[67][30],graph[67][31],graph[67][32],graph[67][33],graph[67][34],graph[67][35],graph[67][36], graph[67][37] , graph[67][38] , graph[67][39] , graph[67][40]  , graph[67][41] , graph[67][42] , graph[67][43] , graph[67][44] , graph[67][45] , graph[67][46] , graph[67][47] , graph[67][48] , graph[67][49] , graph[67][50] , graph[67][51] , graph[67][52] , graph[67][53] , graph[67][54] , graph[67][55] , graph[67][56] , graph[67][57] , graph[67][58] , graph[67][59] , graph[67][60] , graph[67][61] , graph[67][62] , graph[67][63] , graph[67][64] , graph[67][65] , graph[67][66], graph[67][67]} = {6'd60, 6'd60 , 6'd60, 6'd60, 6'd60, 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd60 , 6'd1 , 6'd60 , 6'd60 , 6'd60 , 6'd0};
 end

   
  always@ (posedge clk)
  begin
    if (flag2 != src)
    begin
      dist[0] = 6'd60 ; dist[4] = 6'd60 ; dist[8] = 6'd60 ; dist[12] = 6'd60 ; dist[16] = 6'd60 ; dist[20] = 6'd60 ; dist[24] = 6'd60 ; dist[28] = 6'd60 ; dist[32] = 6'd60 ;
      dist[1] = 6'd60 ; dist[5] = 6'd60 ; dist[9] = 6'd60 ; dist[13] = 6'd60 ; dist[17] = 6'd60 ; dist[21] = 6'd60 ; dist[25] = 6'd60 ; dist[29] = 6'd60 ; dist[33] = 6'd60 ;
      dist[2] = 6'd60 ; dist[6] = 6'd60 ; dist[10] = 6'd60 ; dist[14] = 6'd60 ; dist[18] = 6'd60 ; dist[22] = 6'd60 ; dist[26] = 6'd60 ; dist[30] = 6'd60 ; dist[34] = 6'd60 ;
      dist[3] = 6'd60 ; dist[7] = 6'd60 ; dist[11] = 6'd60 ; dist[15] = 6'd60 ; dist[19] = 6'd60 ; dist[23] = 6'd60 ; dist[27] = 6'd60 ; dist[31] = 6'd60 ; dist[35] = 6'd60 ;
      dist[36] = 6'd60; dist[37] = 6'd60 ; dist[38] = 6'd60 ; dist[39] = 6'd60 ; dist[40] = 6'd60 ; dist[41] = 6'd60 ; dist[42] = 6'd60 ; dist[43] = 6'd60 ; dist[44] = 6'd60 ;
      dist[45] = 6'd60 ; dist[46] = 6'd60 ; dist[47] = 6'd60 ; dist[48] = 6'd60 ; dist[49] = 6'd60 ; dist[50] = 6'd60 ; dist[51] = 6'd60 ; dist[52] = 6'd60 ; dist[53] = 6'd60 ;
      dist[54] = 6'd60 ; dist[55] = 6'd60 ; dist[56] = 6'd60 ; dist[57] = 6'd60 ; dist[58] = 6'd60 ; dist[59] = 6'd60 ; dist[60] = 6'd60 ; dist[61] = 6'd60 ; dist[62] = 6'd60 ;
      dist[63] = 6'd60 ; dist[64] = 6'd60 ; dist[65] = 6'd60 ; dist[66] = 6'd60 ; dist[67] = 6'd60 ;
     
      parent[0] = 7'd60 ; parent[4] = 7'd60 ; parent[8] = 7'd60 ; parent[12] = 7'd60 ; parent[16] = 7'd60 ; parent[20] = 7'd60 ; parent[24] = 7'd60 ; parent[28] = 7'd60 ; parent[32] = 7'd60 ;
      parent[1] = 7'd60 ; parent[5] = 7'd60 ; parent[9] = 7'd60 ; parent[13] = 7'd60 ; parent[17] = 7'd60 ; parent[21] = 7'd60 ; parent[25] = 7'd60 ; parent[29] = 7'd60 ; parent[33] = 7'd60 ;
      parent[2] = 7'd60 ; parent[6] = 7'd60 ; parent[10] = 7'd60 ; parent[14] = 7'd60 ; parent[18] = 7'd60 ; parent[22] = 7'd60 ; parent[26] = 7'd60 ; parent[30] = 7'd60 ; parent[34] = 7'd60 ;
      parent[3] = 7'd60 ; parent[7] = 7'd60 ; parent[11] = 7'd60 ; parent[15] = 7'd60 ; parent[19] = 7'd60 ; parent[23] = 7'd60 ; parent[27] = 7'd60 ; parent[31] = 7'd60 ; parent[35] = 7'd60 ;
      parent[36] = 7'd60; parent[37] = 7'd60 ; parent[38] = 7'd60 ; parent[39] = 7'd60 ; parent[40] = 7'd60 ; parent[41] = 7'd60 ; parent[42] = 7'd60 ; parent[43] = 7'd60 ; parent[44] = 7'd60 ;
      parent[45] = 7'd60 ; parent[46] = 7'd60 ; parent[47] = 7'd60 ; parent[48] = 7'd60 ; parent[49] = 7'd60 ; parent[50] = 7'd60 ; parent[51] = 7'd60 ; parent[52] = 7'd60 ; parent[53] = 7'd60 ;
      parent[54] = 7'd60 ; parent[55] = 7'd60 ; parent[56] = 7'd60 ; parent[57] = 7'd60 ; parent[58] = 7'd60 ; parent[59] = 7'd60 ; parent[60] = 7'd60 ; parent[61] = 7'd60 ; parent[62] = 7'd60 ;
      parent[63] = 7'd60 ; parent[64] = 7'd60 ; parent[65] = 7'd60 ; parent[66] = 7'd60 ; parent[67] = 7'd60 ;

 
      visited = 0 ;
      flag2 = src ;
      path_ready = 0 ;
      path = 0 ;
    end  
    if (temp != src)
    begin
      FindIndex(src,index_src);
      FindIndex(dest,index_dest);
      dist[index_src] = 0 ;
      parent[index_src]= 60 ;  //for our purpose(generally we put -1)
   if (i <= 67 )
   begin
   if(!visited[i] && dist[i]<min)
           begin
            min = dist[i] ;
            key = i ;
           end
   i = i + 1 ;
   end
   if (i > 67)
    begin
      u = key ;
      visited[u] = 1 ;
      if(!visited[v] && (dist[u]+graph[u][v]) <  dist[v] && graph[u][v]!=60)  //60 is infinity in our context
           begin
              parent[v] = u ;
              dist[v] = dist[u] + graph[u][v] ;
           end
       v = v + 1 ;
       if (v == 68)
         begin
          g = g + 1 ;
          v = 0 ;
           i = 0 ;
         key = 0 ;
         min = 60 ;
         end  
       if (g == 67)
         begin
          g = 0 ;
          temp = src ;
          done = 1 ;
          flag = index_dest ;
          j = 1 ;
          //path = 0 ;
         end
    end
    end
    if (done == 1)
    begin
       if (flag == index_dest)
          begin
          temp_index = index_dest ;
          flag = 0 ;
          path[7:0] = dest ;
          end
       if (temp_index != index_src)
       begin
         temp_index = parent[temp_index] ;
         getNode(temp_index,temp_node);
         path[8*j +: 8] = temp_node ;  
         j = j + 1 ;
       end
       else
         begin
         done = 0 ;
         path_ready = 1 ;
         end    
    end
  end

//mapping the nodes
//1-06 2-07 3-08 4-11 5-16 6-17 7-18 8-19 9-22 10-23 11-24 12-26 13-27 14-28 15-30 16-31 17-32 18-33 19-34 20-35 21-42 22-43 23-44 24-52
//25-53 26-54 27-56 28-57 29-58 30-60 31-61 32-62 33-63 34-64 35-65 36-66 37-67 38-68 39-69 40-72 41-73 42-74 43-76 44-77 45-78 46-82 47-83
//48-84 49-90 50-91 51-92 52-93 53-94 54-95 55-102 56-103 57-104 58-106 59-107 60-108 61-111 62-116 63-117 64-118 65-119 66-126 67-127 68-128
//index starts with 0
    task FindIndex ;
    input [7:0] value ;
    output [6:0] index ;
    begin
        case(value[7:4])
                    4'd0 : begin
                              case(value[3:0])
                                 4'd6 : index = 0 ; //06
                                 4'd7 : index = 1 ; //07
                                 4'd8 : index = 2 ; //08
                              endcase
                            end
                     4'd1 : begin
                              case(value[3:0])
                                 4'd1 : index = 3 ; //11
                                 4'd6 : index = 4 ; //16
                                 4'd7 : index = 5 ; //17
                                 4'd8 : index = 6 ; //18
                                 4'd9 : index = 7 ; //19
                              endcase
                            end
                     4'd2 : begin
                              case(value[3:0])
                                 4'd2 : index = 8 ; //22
                                 4'd3 : index = 9 ; //23
                                 4'd4 : index = 10 ; //24
                                 4'd6 : index = 11 ; //26
                                 4'd7 : index = 12 ; //27
                                 4'd8 : index = 13 ; //28
                              endcase
                            end                
                     4'd3 : begin
                              case(value[3:0])
                                 4'd0 : index = 14 ; //30
                                 4'd1 : index = 15 ; //31
                                 4'd2 : index = 16 ; //32
                                 4'd3 : index = 17 ; //33
                                 4'd4 : index = 18 ; //34
                                 4'd5 : index = 19 ; //35
                              endcase
                            end
                     4'd4 : begin
                              case(value[3:0])
                                 4'd2 : index = 20 ; //42
                                 4'd3 : index = 21 ; //43
                                 4'd4 : index = 22 ; //44
                              endcase
                            end    
                     4'd5 : begin
                              case(value[3:0])
                                 4'd2 : index = 23 ; //52
                                 4'd3 : index = 24 ; //53
                                 4'd4 : index = 25 ; //54
                                 4'd6 : index = 26 ; //56
                                 4'd7 : index = 27 ; //57
                                 4'd8 : index = 28 ; //58
                              endcase
                            end            
                     4'd6 : begin
                              case(value[3:0])
                                 4'd0 : index = 29 ; //60
                                 4'd1 : index = 30 ; //61
                                 4'd2 : index = 31 ; //62
                                 4'd3 : index = 32 ; //63
                                 4'd4 : index = 33 ; //64
                                 4'd5 : index = 34 ; //65
                                 4'd6 : index = 35 ; //66
                                 4'd7 : index = 36 ; //67
                                 4'd8 : index = 37 ; //68
                                 4'd9 : index = 38 ; //69
                              endcase
                            end
                      4'd7 : begin
                              case(value[3:0])
                                 4'd2 : index = 39 ; //72
                                 4'd3 : index = 40 ; //73
                                 4'd4 : index = 41 ; //74
                                 4'd6 : index = 42 ; //76
                                 4'd7 : index = 43 ; //77
                                 4'd8 : index = 44 ; //78
                              endcase
                            end
                      4'd8 : begin
                              case(value[3:0])
                                 4'd2 : index = 45 ; //82
                                 4'd3 : index = 46 ; //83
                                 4'd4 : index = 47 ; //84
                              endcase
                            end
                      4'd9 : begin
                              case(value[3:0])
                                 4'd0 : index = 48 ; //90
                                 4'd1 : index = 49 ; //91
                                 4'd2 : index = 50 ; //92
                                 4'd3 : index = 51 ; //93
                                 4'd4 : index = 52 ; //94
                                 4'd5 : index = 53 ; //95
                              endcase
                            end
                      4'd10 : begin
                              case(value[3:0])
                                 4'd2 : index = 54 ; //102
                                 4'd3 : index = 55 ; //103
                                 4'd4 : index = 56 ; //104
                                 4'd6 : index = 57 ; //106
                                 4'd7 : index = 58 ; //107
                                 4'd8 : index = 59 ; //108
                              endcase
end
                      4'd11 : begin
                              case(value[3:0])
                                 4'd1 : index = 60 ; //111
                                 4'd6 : index = 61 ; //116
                                 4'd7 : index = 62 ; //117
                                 4'd8 : index = 63 ; //118
                                 4'd9 : index = 64 ; //119
                              endcase
                            end
                      4'd12 : begin
                              case(value[3:0])
                                 4'd6 : index = 65 ; //126
                                 4'd7 : index = 66 ; //127
                                 4'd8 : index = 67 ; //128
                              endcase
                            end  
endcase
    end
    endtask
   
    task getNode;
     input [6:0] n_index ;
     output [7:0] node ;
     begin
      case(n_index)
        7'd0 : node = {4'd0,4'd6} ; //06
        7'd1 : node = {4'd0,4'd7} ; //07
        7'd2 : node = {4'd0,4'd8} ; //08
        7'd3 : node = {4'd1,4'd1} ; //11
        7'd4 : node = {4'd1,4'd6} ; //16
        7'd5 : node = {4'd1,4'd7} ; //17
        7'd6 : node = {4'd1,4'd8} ; //18
        7'd7 : node = {4'd1,4'd9} ; //19
        7'd8 : node = {4'd2,4'd2} ; //22
        7'd9 : node = {4'd2,4'd3} ; //23
        7'd10 : node = {4'd2,4'd4} ; //24
        7'd11 : node = {4'd2,4'd6} ; //26
        7'd12 : node = {4'd2,4'd7} ; //27
        7'd13 : node = {4'd2,4'd8} ; //28
        7'd14 : node = {4'd3,4'd0} ; //30
        7'd15 : node = {4'd3,4'd1} ; //31
        7'd16 : node = {4'd3,4'd2} ; //32
        7'd17 : node = {4'd3,4'd3} ; //33
        7'd18 : node = {4'd3,4'd4} ; //34
        7'd19 : node = {4'd3,4'd5} ; //35
        7'd20 : node = {4'd4,4'd2} ; //42
        7'd21 : node = {4'd4,4'd3} ; //43
        7'd22 : node = {4'd4,4'd4} ; //44
        7'd23 : node = {4'd5,4'd2} ; //52
        7'd24 : node = {4'd5,4'd3} ; //53
        7'd25 : node = {4'd5,4'd4} ; //54
        7'd26 : node = {4'd5,4'd6} ; //56
        7'd27 : node = {4'd5,4'd7} ; //57
        7'd28 : node = {4'd5,4'd8} ; //58
        7'd29 : node = {4'd6,4'd0} ; //60
        7'd30 : node = {4'd6,4'd1} ; //61
        7'd31 : node = {4'd6,4'd2} ; //62
        7'd32 : node = {4'd6,4'd3} ; //63
        7'd33 : node = {4'd6,4'd4} ; //64
        7'd34 : node = {4'd6,4'd5} ; //65
        7'd35 : node = {4'd6,4'd6} ; //66
        7'd36 : node = {4'd6,4'd7} ; //67
        7'd37 : node = {4'd6,4'd8} ; //68
        7'd38 : node = {4'd6,4'd9} ; //69
        7'd39 : node = {4'd7,4'd2} ; //72
        7'd40 : node = {4'd7,4'd3} ; //73
        7'd41 : node = {4'd7,4'd4} ; //74
        7'd42 : node = {4'd7,4'd6} ; //76
        7'd43 : node = {4'd7,4'd7} ; //77
        7'd44 : node = {4'd7,4'd8} ; //78
        7'd45 : node = {4'd8,4'd2} ; //82
        7'd46 : node = {4'd8,4'd3} ; //83
        7'd47 : node = {4'd8,4'd4} ; //84
        7'd48 : node = {4'd9,4'd0} ; //90
        7'd49 : node = {4'd9,4'd1} ; //91
        7'd50 : node = {4'd9,4'd2} ; //92
        7'd51 : node = {4'd9,4'd3} ; //93
        7'd52 : node = {4'd9,4'd4} ; //94
        7'd53 : node = {4'd9,4'd5} ; //95
        7'd54 : node = {4'd10,4'd2} ; //102
        7'd55 : node = {4'd10,4'd3} ; //103
        7'd56 : node = {4'd10,4'd4} ; //104
        7'd57 : node = {4'd10,4'd5} ; //105
        7'd58 : node = {4'd10,4'd7} ; //107
        7'd59 : node = {4'd10,4'd8} ; //108
        7'd60 : node = {4'd11,4'd1} ; //111
        7'd61 : node = {4'd11,4'd6} ; //116
        7'd62 : node = {4'd11,4'd7} ; //117
        7'd63 : node = {4'd11,4'd8} ; //118
        7'd64 : node = {4'd11,4'd9} ; //119
        7'd65 : node = {4'd12,4'd6} ; //126
        7'd66 : node = {4'd12,4'd7} ; //127
        7'd67 : node = {4'd12,4'd8} ; //128
      endcase
     end
    endtask

   
endmodule
